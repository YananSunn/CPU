`timescale 1ns / 1ps

module vga
#(parameter WIDTH = 0, HSIZE = 800, HFP = 856, HSP = 976, HMAX = 1040, VSIZE = 600, VFP = 637, VSP = 643, VMAX = 666, HSPP = 1, VSPP = 1)
(
    input wire clk,
    input wire enable,
    input wire[19199:0] signal_input,
    input wire[31:0] char_pos,
    output wire[2:0] video_red,    
    output wire[2:0] video_green,  
    output wire[1:0] video_blue,   
    output wire video_hsync,       
    output wire video_vsync,       
    output wire video_clk,         
    output wire video_de           
);
    reg [11:0] hdata;
    reg [11:0] vdata;
    reg [6:0] flag;
    reg [6:0] hpos;
    reg [6:0] vpos;
    reg [6:0] hcount;
    reg [6:0] vcount;
    assign video_clk = clk;
    reg [199:0] character;

    reg hof_flag,vof_flag;

    reg[2:0] videored;   
    reg[2:0] videogreen; 
    reg[1:0] videoblue;  
    wire[7:0] char_index;
    assign char_index[0] = signal_input[vpos * 640 + hpos * 8];
    assign char_index[1] = signal_input[vpos * 640 + hpos * 8 + 1];
    assign char_index[2] = signal_input[vpos * 640 + hpos * 8 + 2];
    assign char_index[3] = signal_input[vpos * 640 + hpos * 8 + 3];
    assign char_index[4] = signal_input[vpos * 640 + hpos * 8 + 4];
    assign char_index[5] = signal_input[vpos * 640 + hpos * 8 + 5];
    assign char_index[6] = signal_input[vpos * 640 + hpos * 8 + 6];
    assign char_index[7] = signal_input[vpos * 640 + hpos * 8 + 7];
    always @(posedge clk) begin
        if(enable)begin
            if(vof_flag || hof_flag)begin
                videored <= 3'b000;
                videogreen <= 3'b000;
                videoblue <= 2'b00;
            end
            else begin
                case (char_index)
                    8'b00100001:
                            character <= 200'b11111111111111111111111111111111111111111111001111111100111111111111111111001111111100111111110011111110000111111000011111100001111110000111111000011111110011111111111111111111111111111111111111111111 ;
					8'b00100010:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011110011001111001100111111111111111111111111111111111111111111 ;
					8'b00100011:
							character <= 200'b11111111111111111111111111111111111111111100110011110011001111001100111000000001100000000111001100111100110011100000000110000000011100110011110011001111001100111111111111111111111111111111111111111111 ;
					8'b00100100:
							character <= 200'b11111111111111111111111100111111110011111110000111110000001110001100011000111111110011111111100111111111000111111110001111111100011000110001110000001111100001111111001111111100111111111111111111111111 ;
					8'b00100101:
							character <= 200'b11111111111111111111111111111111111111111000111001001001100100001100111000110011111110000111111001111111001111111100111111100111111110010001110010010011001001001111110001111111111111111111111111111111 ;
					8'b00100110:
							character <= 200'b11111111111111111111111111111111111111110010000111100000001111001110011101111001100111100100001100111111100111111000111111001001111001110011110010011111100011111111111111111111111111111111111111111111 ;
					8'b00100111:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100111111110011111111111111111111111111111111111111111111 ;
					8'b00101000:
							character <= 200'b11111111111110011111111100111111111001111111110111111111001111111100111111110011111111001111111100111111110011111111001111111100111111110111111110011111110011111110011111111111111111111111111111111111 ;
					8'b00101001:
							character <= 200'b11111111111111110011111110011111110011111111011111111001111111100111111110011111111001111111100111111110011111111001111111100111111111011111111100111111111001111111110011111111111111111111111111111111 ;
					8'b00101010:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111110011110011100110011111000011110000000011110000111110011001110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00101011:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111001111111100111111110011111000000001100000000111110011111111001111111100111111111111111111111111111111111111111111111111111111 ;
					8'b00101100:
							character <= 200'b11111111111111111111111110111111110111111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00101101:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00101110:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00101111:
							character <= 200'b11111111111111111111111111100111111110011111110011111111001111111001111111100111111100111111110011111110011111111001111111001111111100111111100111111110011111111111111111111111111111111111111111111111 ;
					8'b00110000:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100111100110010010011001001001100111100110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00110001:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111000011111100001111110011111111111111111111111111111111111111111111 ;
					8'b00110010:
							character <= 200'b11111111111111111111111111111111111111111000000001100000000111111100011111100011111100011111100011111100011111100011111110011111111000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00110011:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111111100011111111000011111110001111110011111110011111111000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00110100:
							character <= 200'b11111111111111111111111111111111111111111100111111110011111111001111111100111111100000000110000000011100111001110011001111001100111100110011110011001111111100111111111111111111111111111111111111111111 ;
					8'b00110101:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111111100111111110001111111100000001111000000111111110011111111001100000000110000000011111111111111111111111111111111111111111 ;
					8'b00110110:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100011000111000000011110001001111111100111111110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00110111:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111110011111111001111111100111111110011111111001111111001111111001111111001111111100000001110000000111111111111111111111111111111111111111111 ;
					8'b00111000:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100011000111000000111110000111110011001110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00111001:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111111100111111110001001111000000011100011000110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b00111010:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111111111111111111111111111111111110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00111011:
							character <= 200'b11111111111111111111111110111111110111111111001111111100111111111111111111111111111111111111110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00111100:
							character <= 200'b11111111111111111111111111111111111111111100111111111001111111110011111111100111111111001111111110011111110011111110011111110011111110011111110011111111111111111111111111111111111111111111111111111111 ;
					8'b00111101:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111110000011111000001111111111111111111111111000001111100000111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b00111110:
							character <= 200'b11111111111111111111111111111111111111111111110011111110011111110011111110011111110011111110011111111100111111111001111111110011111111100111111111001111111111111111111111111111111111111111111111111111 ;
					8'b00111111:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111111111111111001111111100111111100011111100011111100011111110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01000000:
							character <= 200'b11111111111111111111111111111110000001111000000011111111100110000110011000001001100110100110011010011000001001100001100110011110011001111001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01000001:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011000000001100000000110011110011001111001100111100110011110011100110011111000011111110011111111111111111111111111111111111111111111 ;
					8'b01000010:
							character <= 200'b11111111111111111111111111111111111111111110000001110000000110011110011001111001100111100111000000011100000001100111100110011110011001111001110000000111100000011111111111111111111111111111111111111111 ;
					8'b01000011:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011111111001111111100111111110011111111001111111100111111110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01000100:
							character <= 200'b11111111111111111111111111111111111111111110000001110000000110001110011001111001100111100110011110011001111001100111100110011110011000111001110000000111100000011111111111111111111111111111111111111111 ;
					8'b01000101:
							character <= 200'b11111111111111111111111111111111111111111000000001100000000111111110011111111001111111100111100000011110000001111111100111111110011111111001100000000110000000011111111111111111111111111111111111111111 ;
					8'b01000110:
							character <= 200'b11111111111111111111111111111111111111111111111001111111100111111110011111111001111111100111100000011110000001111111100111111110011111111001100000000110000000011111111111111111111111111111111111111111 ;
					8'b01000111:
							character <= 200'b11111111111111111111111111111111111111111001000111100000001110001100011001111001100001100110000110011111111001111111100111111110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01001000:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011001111001100111100110000000011000000001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01001001:
							character <= 200'b11111111111111111111111111111111111111111100000011110000001111110011111111001111111100111111110011111111001111111100111111110011111111001111110000001111000000111111111111111111111111111111111111111111 ;
					8'b01001010:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111111111111111111111111111111111111111111 ;
					8'b01001011:
							character <= 200'b11111111111111111111111111111111111111111001111001100011100111000110011110001001111100000111111000011111110001111110000111110000011110001001110001100111001110011111111111111111111111111111111111111111 ;
					8'b01001100:
							character <= 200'b11111111111111111111111111111111111111111000000001100000000111111110011111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111111111111111111111111111111111111 ;
					8'b01001101:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011001111001100100100110010010011000000001100000000110001100011000110001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01001110:
							character <= 200'b11111111111111111111111111111111111111111001111001100011100110001110011000011001100001100110010010011001001001100110000110011000011001110001100111000110011110011111111111111111111111111111111111111111 ;
					8'b01001111:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100111100110011110011001111001100111100110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01010000:
							character <= 200'b11111111111111111111111111111111111111111111111001111111100111111110011111111001111000000111000000011000111001100111100110011110011000111001110000000111100000011111111111111111111111111111111111111111 ;
					8'b01010001:
							character <= 200'b11111111111111111111111111111111111111111001000111100000001110000100011000011001100111100110011110011001111001100111100110011110011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01010010:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011100111001111000000111000000011000111001100111100110011110011000111001110000000111100000011111111111111111111111111111111111111111 ;
					8'b01010011:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011000111111110011111111100111111111000111111110001111111100011000110001110000001111100001111111111111111111111111111111111111111111 ;
					8'b01010100:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111001111100000000110000000011111111111111111111111111111111111111111 ;
					8'b01010101:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100111100110011110011001111001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01010110:
							character <= 200'b11111111111111111111111111111111111111111111001111111000011111001100111001111001100111100110011110011001111001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01010111:
							character <= 200'b11111111111111111111111111111111111111111100110011100000000110010010011001001001100100100110010010011001001001100100100110011110011001111001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01011000:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100111001100111100110011111000011111110011111111001111111000011111001100111100110011100111100110011110011111111111111111111111111111111111111111 ;
					8'b01011001:
							character <= 200'b11111111111111111111111111111111111111111111001111111100111111110011111111001111111100111111100001111100110011100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111 ;
					8'b01011010:
							character <= 200'b11111111111111111111111111111111111111111000000001100000000111111110011111110001111110001111110001111110001111110001111110001111111001111111100000000110000000011111111111111111111111111111111111111111 ;
					8'b01011011:
							character <= 200'b11111111111110000111111000011111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111001111111100111111000011111100001111111111111111111111111111111111111111111 ;
					8'b01011100:
							character <= 200'b11111111111111111111100111111110011111111100111111110011111111100111111110011111111100111111110011111111100111111110011111111100111111110011111111100111111110011111111111111111111111111111111111111111 ;
					8'b01011101:
							character <= 200'b11111111111110000111111000011111100111111110011111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111000011111100001111111111111111111111111111111111111111111 ;
					8'b01011110:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011100110011111000011111110011111111111111 ;
					8'b01011111:
							character <= 200'b11111111111000000001100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01100000:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100111111110001111111111111 ;
					8'b01100001:
							character <= 200'b11111111111111111111111111111111111111111000000011100000000110011110011001111001100000000110000000111001111111110000001111100000111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01100010:
							character <= 200'b11111111111111111111111111111111111111111110001001110000000110001100011001111001100111100110011110011000110001110000000111100010011111111001111111100111111110011111111111111111111111111111111111111111 ;
					8'b01100011:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011111111001111111100111111110011000110001110000001111100001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01100100:
							character <= 200'b11111111111111111111111111111111111111111001000111100000001110001100011001111001100111100110011110011000110001100000001110010001111001111111100111111110011111111111111111111111111111111111111111111111 ;
					8'b01100101:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001111111100011000000001100000000110011110011000110001110000001111100001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01100110:
							character <= 200'b11111111111111111111111111111111111111111111100111111110011111111001111111100111111110011111111001111000000001100000000111111001111111100111100000011110000011111111111111111111111111111111111111111111 ;
					8'b01100111:
							character <= 200'b11100000111100000011100011111110011111111001000111100000001110001100011001111001100111100110011110011000110001110000001111100001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01101000:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011001111001100111100110011110011000110001110000000111100010011111111001111111100111111110011111111111111111111111111111111111111111 ;
					8'b01101001:
							character <= 200'b11111111111111111111111111111111111111111100000011110000001111110011111111001111111100111111110011111111001111111100001111110000111111111111111111111111110011111111001111111111111111111111111111111111 ;
					8'b01101010:
							character <= 200'b11111000111111000011111000111111100111111110011111111001111111100111111110011111111001111111100111111110011111111000011111100001111111111111111111111111100111111110011111111111111111111111111111111111 ;
					8'b01101011:
							character <= 200'b11111111111111111111111111111111111111111001111001110011100111100110011111000001111111000111111000011111001001111001100111001110011111111001111111100111111110011111111111111111111111111111111111111111 ;
					8'b01101100:
							character <= 200'b11111111111111111111111111111111111111111100000011110000001111110011111111001111111100111111110011111111001111111100111111110011111111001111111100001111110000111111111111111111111111111111111111111111 ;
					8'b01101101:
							character <= 200'b11111111111111111111111111111111111111111001001001100100100110010010011001001001100100100110010010011001001001100000000111010010011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01101110:
							character <= 200'b11111111111111111111111111111111111111111001111001100111100110011110011001111001100111100110011110011000110001110000000111100010011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01101111:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110001100011001111001100111100110011110011000110001110000001111100001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110000:
							character <= 200'b11111110011111111001111111100111111110011110001001110000000110001100011001111001100111100110011110011000110001110000000111100010011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110001:
							character <= 200'b10011111111001111111100111111110011111111001000111100000001110001100011001111001100111100110011110011000110001100000001110010001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110010:
							character <= 200'b11111111111111111111111111111111111111111111111001111111100111111110011111111001111111100111111100011111100001100000000110000010011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110011:
							character <= 200'b11111111111111111111111111111111111111111110000111110000001110011110011000111111110000001111111100011001111001110000001111100001111111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110100:
							character <= 200'b11111111111111111111111111111111111111111100001111110000011111111001111111100111111110011111111001111111100111110000001111000000111111100111111110011111111001111111111111111111111111111111111111111111 ;
					8'b01110101:
							character <= 200'b11111111111111111111111111111111111111111001000111100000001110001100011001111001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110110:
							character <= 200'b11111111111111111111111111111111110011111110000111110011001110011110011001111001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01110111:
							character <= 200'b11111111111111111111111111111111111111111101111011100011000110000000011000000001100100100110010010011001111001100111100110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01111000:
							character <= 200'b11111111111111111111111111111111111111111001111001100011000111000000111110000111111100111111100001111100000011100011000110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01111001:
							character <= 200'b11100000111100000011100111111110011111111001000111100000001110001100011001111001100111100110011110011001111001100111100110011110011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01111010:
							character <= 200'b11111111111111111111111111111111111111111000000001100000000111111100111111100111111100111111100111111100111111100000000110000000011111111111111111111111111111111111111111111111111111111111111111111111 ;
					8'b01111011:
							character <= 200'b11111111111100011111111100111111111001111111100111111110011111111001111111100111111111001111111001111111100111111110011111111001111111100111111100111111000111111111111111111111111111111111111111111111 ;
					8'b01111100:
							character <= 200'b11111111111111111111111111111111110011111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111001111111100111111110011111111111111111111111111111111111111111111 ;
					8'b01111101:
							character <= 200'b11111111111111100011111100111111100111111110011111111001111111100111111110011111110011111111100111111110011111111001111111100111111110011111111100111111111000111111111111111111111111111111111111111111 ;
					8'b01111110:
							character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011101100100100110111000111111111111111111111111111111111111111111 ;
					default:
						character <= 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 ;
                endcase
                if((hpos == char_pos[22:16]) && (vpos == char_pos[6:0]) && (hcount < 3))begin
                    if(character[vcount*10+hcount] == 1)begin
                        videored <= 3'b000;
                        videogreen <= 3'b000;
                        videoblue <= 2'b00;
                    end
                    else begin
                        videored <= 3'b111;
                        videogreen <= 3'b111;
                        videoblue <= 2'b11;
                    end
                end
                else begin
                    if(character[vcount*10+hcount] == 1)begin
                        videored <= 3'b111;
                        videogreen <= 3'b111;
                        videoblue <= 2'b11;
                    end
                    else begin
                        videored <= 3'b000;
                        videogreen <= 3'b000;
                        videoblue <= 2'b00;
                    end
                end
            end
        end
    end

    // init
    initial begin
        hdata <= 0;
        vdata <= 0;
        hpos <= 0;
        vpos <= 0;
        hcount <= 0;
        vcount <= 0;
    end

    // hdata
    always @ (posedge clk)
    begin
        if (hdata >= (HMAX - 1))begin
            hdata <= 0;
        end
        else begin
            hdata <= hdata + 1;
        end
        if(hdata < 800)begin
            hof_flag <= 0;
            if (hcount >= 9) begin
                hcount <= 0;
                if (hpos >= 79)
                    hpos <= 0;
                else
                    hpos <= hpos + 1;
            end
            else begin
                hcount <= hcount+1;
            end
        end
        else begin
            hof_flag <= 1;
        end
    end

    // vdata
    always @ (posedge clk)
    begin
        if (hdata >= (HMAX - 1)) 
        begin
            if (vdata >= (VMAX - 1))begin
                vdata <= 0;
            end
            else begin
                vdata <= vdata + 1;
            end

            if(vdata < 600)begin
                vof_flag <= 0;
                if (vcount >= 19) begin
                    vcount <= 0;
                    if (vpos >= 29)
                        vpos <= 0;
                    else
                        vpos <= vpos + 1;
                end
                else begin
                    vcount <= vcount+1;
                end
            end
            else begin
                vof_flag <= 1;
            end
        end
    end

    // hsync & vsync & blank
    assign video_hsync = ((hdata >= HFP) && (hdata < HSP)) ? HSPP : !HSPP;
    assign video_vsync = ((vdata >= VFP) && (vdata < VSP)) ? VSPP : !VSPP;
    assign video_de = ((hdata < HSIZE) & (vdata < VSIZE));
    assign video_red    = videored;
    assign video_green  = videogreen;
    assign video_blue   = videoblue;

endmodule