module MMU(
    input wire clk,
    
    input wire if_read,
    input wire if_write,
    input wire[31:0] addr,
    input wire[31:0] input_data,
    input wire bytemode,
    output reg[31:0] output_data,
    
    inout wire[31:0] base_ram_data,
    output wire[19:0] base_ram_addr,
    output wire[3:0] base_ram_be_n,
    output wire base_ram_ce_n,
    output wire base_ram_oe_n,
    output wire base_ram_we_n,

    inout wire[31:0] ext_ram_data,
    output wire[19:0] ext_ram_addr,
    output wire[3:0] ext_ram_be_n,
    output wire ext_ram_ce_n,
    output wire ext_ram_oe_n,
    output wire ext_ram_we_n,
    
    output wire uart_rdn,
    output wire uart_wrn,
    input wire uart_dataready,
    input wire uart_tbre,
    input wire uart_tsre
    );

reg oe1 = 1'b1, we1 = 1'b1, ce1 = 1'b1;
reg oe2 = 1'b1, we2 = 1'b1, ce2 = 1'b1;
reg[3:0] be = 4'b0000;
reg[31:0] ram_read_data1, ram_read_data2, ram_write_data;
reg wrn = 1'b1, rdn = 1'b1;

assign base_ram_addr = addr[21:2];
assign ext_ram_addr  = addr[21:2];

assign base_ram_data = if_write ? ram_write_data :  32'bz;
assign ext_ram_data  = if_write ? ram_write_data :  32'bz;

assign base_ram_ce_n = ce1;
assign base_ram_oe_n = oe1;
assign base_ram_we_n = we1;
assign base_ram_be_n = be;

assign ext_ram_ce_n = ce2;
assign ext_ram_oe_n = oe2;
assign ext_ram_we_n = we2;
assign ext_ram_be_n = be;

assign uart_wrn     = wrn;
assign uart_rdn     = rdn;

wire[31:0] ram_read_data = addr[22] ? ext_ram_data : base_ram_data;

always @(*) begin
    if (clk) begin
        case (addr)
            32'hBFD003F8: begin
                ce1 <= 1'b1;
                ce2 <= 1'b1;
                if (if_read) begin
                    rdn <= 1'b0;
                    wrn <= 1'b1;
                    output_data <= {24'b0, base_ram_data[7:0]};
                end
                else if (if_write) begin
                    rdn <= 1'b1;
                    wrn <= 1'b0;
                    ram_write_data <= input_data;
                end
                else begin
                    rdn <= 1'b1;
                    wrn <= 1'b1;
                end
            end
            32'hBFD003FD: begin
                ce1 <= 1'b1;
                ce2 <= 1'b1;
                rdn <= 1'b1;
                wrn <= 1'b1;
                if (if_read) begin
                    output_data <= {30'b0, uart_dataready, uart_tsre};
                end
            end
            default: begin
                // RAM
                ce1 <= addr[22];
                ce2 <= ~addr[22];
                oe1 <= addr[22] | (~if_read);
                oe2 <= (~addr[22]) | (~if_read);
                we1 <= addr[22] | (~if_write);
                we2 <= (~addr[22]) | (~if_write);
                rdn <= 1'b1;
                wrn <= 1'b1;
                if (if_read) begin
                    if (bytemode) begin
                        case (addr[1:0])
                            2'b00: begin
                                output_data <= {{24{ram_read_data[31]}}, ram_read_data[31:24]};
                                be <= 4'b0111;
                            end
                            2'b01: begin
                                output_data <= {{24{ram_read_data[23]}}, ram_read_data[23:16]};
                                be <= 4'b1011;
                            end
                            2'b10: begin
                                output_data <= {{24{ram_read_data[15]}}, ram_read_data[15:8]};
                                be <= 4'b1101;
                            end
                            2'b11: begin
                                output_data <= {{24{ram_read_data[7]}}, ram_read_data[7:0]};
                                be <= 4'b1110;
                            end
                            default: begin
                                output_data <= ram_read_data;
                                be <= 4'b0000;
                            end
                        endcase
                    end
                    else begin
/*
                    // for DEBUG
                        case (addr)
                            32'h80000000: output_data <= 32'b00111100000110101000000000000000;
                            32'h80000004: output_data <= 32'b00100111010110100001000110111100;
                            32'h80000008: output_data <= 32'b00000011010000000000000000001000;
                            32'h80001180: output_data <= 32'b00111100000110101000000000000000;
                            32'h80001184: output_data <= 32'b00100111010110100001010111000100;
                            32'h80001188: output_data <= 32'b00000011010000000000000000001000;
                            32'h80001190: output_data <= 32'b01001001010011100100111101001101;
                            32'h80001194: output_data <= 32'b00100000010100100100111101010100;
                            32'h80001198: output_data <= 32'b00100000011100100110111101100110;
                            32'h8000119C: output_data <= 32'b01010011010100000100100101001101;
                            32'h800011A0: output_data <= 32'b00101101001000000011001000110011;
                            32'h800011A4: output_data <= 32'b01101001011011100110100100100000;
                            32'h800011A8: output_data <= 32'b01101100011000010110100101110100;
                            32'h800011AC: output_data <= 32'b01100100011001010111101001101001;
                            32'h800011B0: output_data <= 32'b00000000000000000000000000101110;
                            32'h800011B4: output_data <= 32'b10000000011111110000000000000000;
                            32'h800011B8: output_data <= 32'b10000000011111110000000010001100;
                            32'h800011BC: output_data <= 32'b00111100000110101000000001111111;
                            32'h800011C0: output_data <= 32'b00100111010110100000000000000000;
                            32'h800011C4: output_data <= 32'b00111100000110111000000001111111;
                            32'h800011C8: output_data <= 32'b00100111011110110000000010001100;
                            32'h800011CC: output_data <= 32'b00010011010110110000000000000101;
                            32'h800011D4: output_data <= 32'b10101111010000000000000000000000;
                            32'h800011D8: output_data <= 32'b00100111010110100000000000000100;
                            32'h800011DC: output_data <= 32'b00010000000000001111111111111011;
                            32'h800011E4: output_data <= 32'b00111100000111011000000010000000;
                            32'h800011E8: output_data <= 32'b00100111101111010000000000000000;
                            32'h800011EC: output_data <= 32'b00000011101000001111000000100101;
                            32'h800011F0: output_data <= 32'b00111100000010001000000001111111;
                            32'h800011F4: output_data <= 32'b00100101000010000000000000000000;
                            32'h800011F8: output_data <= 32'b00111100000010011000000001111111;
                            32'h800011FC: output_data <= 32'b10101101001010000000000001110000;
                            32'h80001200: output_data <= 32'b00111100000010011000000001111111;
                            32'h80001204: output_data <= 32'b10101101001010000000000001110100;
                            32'h80001208: output_data <= 32'b00111100000010001011111111010000;
                            32'h8000120C: output_data <= 32'b00110100000010010000000000010000;
                            32'h80001210: output_data <= 32'b10100001000010010000001111111100;
                            32'h80001214: output_data <= 32'b00110100000010000000000000100000;
                            32'h80001218: output_data <= 32'b00100101000010001111111111111111;
                            32'h8000121C: output_data <= 32'b00100111101111011111111111111100;
                            32'h80001220: output_data <= 32'b10101111101000000000000000000000;
                            32'h80001224: output_data <= 32'b00010101000000001111111111111100;
                            32'h8000122C: output_data <= 32'b00111100000010001000000001111111;
                            32'h80001230: output_data <= 32'b00100101000010000000000010000000;
                            32'h80001234: output_data <= 32'b10101101000111010000000000000000;
                            32'h80001238: output_data <= 32'b00000011101000000111000000100101;
                            32'h8000123C: output_data <= 32'b00110100000010000000000000100000;
                            32'h80001240: output_data <= 32'b00100101000010001111111111111111;
                            32'h80001244: output_data <= 32'b00100111101111011111111111111100;
                            32'h80001248: output_data <= 32'b10101111101000000000000000000000;
                            32'h8000124C: output_data <= 32'b00010101000000001111111111111100;
                            32'h80001254: output_data <= 32'b00111100000010001000000001111111;
                            32'h80001258: output_data <= 32'b00100101000010000000000010000000;
                            32'h8000125C: output_data <= 32'b10101101000111010000000000000100;
                            32'h80001260: output_data <= 32'b10101101110111010000000001111100;
                            32'h80001264: output_data <= 32'b00111100000010101000000001111111;
                            32'h80001268: output_data <= 32'b00100101010010100000000010000100;
                            32'h8000126C: output_data <= 32'b10001101010010100000000000000000;
                            32'h80001270: output_data <= 32'b00111100000010011000000001111111;
                            32'h80001274: output_data <= 32'b10101101001010100000000010001000;
                            32'h80001278: output_data <= 32'b00001000000000000000010010100000;
                            32'h80001280: output_data <= 32'b00111100000100001000000000000000;
                            32'h80001284: output_data <= 32'b00100110000100000001000110010000;
                            32'h80001288: output_data <= 32'b10000010000001000000000000000000;
                            32'h8000128C: output_data <= 32'b00100110000100000000000000000001;
                            32'h80001290: output_data <= 32'b00001100000000000000010101110011;
                            32'h80001298: output_data <= 32'b10000010000001000000000000000000;
                            32'h8000129C: output_data <= 32'b00010100100000001111111111111011;
                            32'h800012A4: output_data <= 32'b00001000000000000000010010111001;
                            32'h800012D4: output_data <= 32'b00001000000000000000010010101011;
                            32'h800012DC: output_data <= 32'b00010000000000001111111111111111;
                            32'h800012E4: output_data <= 32'b00001100000000000000010101111110;
                            32'h800012EC: output_data <= 32'b00110100000010000000000001010010;
                            32'h800012F0: output_data <= 32'b00010000010010000000000000100110;
                            32'h800012F8: output_data <= 32'b00110100000010000000000001000100;
                            32'h800012FC: output_data <= 32'b00010000010010000000000000110100;
                            32'h80001304: output_data <= 32'b00110100000010000000000001000001;
                            32'h80001308: output_data <= 32'b00010000010010000000000001000110;
                            32'h80001310: output_data <= 32'b00110100000010000000000001000111;
                            32'h80001314: output_data <= 32'b00010000010010000000000001011001;
                            32'h8000131C: output_data <= 32'b00110100000010000000000001010100;
                            32'h80001320: output_data <= 32'b00010000010010000000000000000011;
                            32'h80001328: output_data <= 32'b00001000000000000000010101101111;
                            32'h80001330: output_data <= 32'b00001100000000000000010110001001;
                            32'h80001338: output_data <= 32'b00100111101111011111111111101000;
                            32'h8000133C: output_data <= 32'b10101111101100000000000000000000;
                            32'h80001340: output_data <= 32'b10101111101100010000000000000100;
                            32'h80001344: output_data <= 32'b00100100000100001111111111111111;
                            32'h80001348: output_data <= 32'b10101111101100000000000000001100;
                            32'h8000134C: output_data <= 32'b10101111101100000000000000010000;
                            32'h80001350: output_data <= 32'b10101111101100000000000000010100;
                            32'h80001354: output_data <= 32'b00110100000100010000000000001100;
                            32'h80001358: output_data <= 32'b00100111101100000000000000001100;
                            32'h8000135C: output_data <= 32'b10000010000001000000000000000000;
                            32'h80001360: output_data <= 32'b00100110001100011111111111111111;
                            32'h80001364: output_data <= 32'b00001100000000000000010101110011;
                            32'h8000136C: output_data <= 32'b00100110000100000000000000000001;
                            32'h80001370: output_data <= 32'b00010110001000001111111111111010;
                            32'h80001378: output_data <= 32'b10001111101100000000000000000000;
                            32'h8000137C: output_data <= 32'b10001111101100010000000000000100;
                            32'h80001380: output_data <= 32'b00100111101111010000000000011000;
                            32'h80001384: output_data <= 32'b00001000000000000000010101101111;
                            32'h8000138C: output_data <= 32'b00100111101111011111111111111000;
                            32'h80001390: output_data <= 32'b10101111101100000000000000000000;
                            32'h80001394: output_data <= 32'b10101111101100010000000000000100;
                            32'h80001398: output_data <= 32'b00111100000100001000000001111111;
                            32'h8000139C: output_data <= 32'b00110100000100010000000001111000;
                            32'h800013A0: output_data <= 32'b10000010000001000000000000000000;
                            32'h800013A4: output_data <= 32'b00100110001100011111111111111111;
                            32'h800013A8: output_data <= 32'b00001100000000000000010101110011;
                            32'h800013B0: output_data <= 32'b00100110000100000000000000000001;
                            32'h800013B4: output_data <= 32'b00010110001000001111111111111010;
                            32'h800013BC: output_data <= 32'b10001111101100000000000000000000;
                            32'h800013C0: output_data <= 32'b10001111101100010000000000000100;
                            32'h800013C4: output_data <= 32'b00100111101111010000000000001000;
                            32'h800013C8: output_data <= 32'b00001000000000000000010101101111;
                            32'h800013D0: output_data <= 32'b00100111101111011111111111111000;
                            32'h800013D4: output_data <= 32'b10101111101100000000000000000000;
                            32'h800013D8: output_data <= 32'b10101111101100010000000000000100;
                            32'h800013DC: output_data <= 32'b00001100000000000000010110001001;
                            32'h800013E4: output_data <= 32'b00000000010000001000000000100101;
                            32'h800013E8: output_data <= 32'b00001100000000000000010110001001;
                            32'h800013F0: output_data <= 32'b00000000010000001000100000100101;
                            32'h800013F4: output_data <= 32'b10000010000001000000000000000000;
                            32'h800013F8: output_data <= 32'b00100110001100011111111111111111;
                            32'h800013FC: output_data <= 32'b00001100000000000000010101110011;
                            32'h80001404: output_data <= 32'b00100110000100000000000000000001;
                            32'h80001408: output_data <= 32'b00010110001000001111111111111010;
                            32'h80001410: output_data <= 32'b10001111101100000000000000000000;
                            32'h80001414: output_data <= 32'b10001111101100010000000000000100;
                            32'h80001418: output_data <= 32'b00100111101111010000000000001000;
                            32'h8000141C: output_data <= 32'b00001000000000000000010101101111;
                            32'h80001424: output_data <= 32'b00100111101111011111111111111000;
                            32'h80001428: output_data <= 32'b10101111101100000000000000000000;
                            32'h8000142C: output_data <= 32'b10101111101100010000000000000100;
                            32'h80001430: output_data <= 32'b00001100000000000000010110001001;
                            32'h80001438: output_data <= 32'b00000000010000001000000000100101;
                            32'h8000143C: output_data <= 32'b00001100000000000000010110001001;
                            32'h80001444: output_data <= 32'b00000000010000001000100000100101;
                            32'h80001448: output_data <= 32'b00000000000100011000100010000010;
                            32'h8000144C: output_data <= 32'b00001100000000000000010110001001;
                            32'h80001454: output_data <= 32'b10101110000000100000000000000000;
                            32'h80001458: output_data <= 32'b00100110001100011111111111111111;
                            32'h8000145C: output_data <= 32'b00100110000100000000000000000100;
                            32'h80001460: output_data <= 32'b00010110001000001111111111111010;
                            32'h80001468: output_data <= 32'b10001111101100000000000000000000;
                            32'h8000146C: output_data <= 32'b10001111101100010000000000000100;
                            32'h80001470: output_data <= 32'b00100111101111010000000000001000;
                            32'h80001474: output_data <= 32'b00001000000000000000010101101111;
                            32'h8000147C: output_data <= 32'b00001100000000000000010110001001;
                            32'h80001484: output_data <= 32'b00110100000001000000000000000110;
                            32'h80001488: output_data <= 32'b00001100000000000000010101110011;
                            32'h80001490: output_data <= 32'b00000000010000001101000000100101;
                            32'h80001494: output_data <= 32'b00111100000111111000000001111111;
                            32'h80001498: output_data <= 32'b00100111111111110000000000000000;
                            32'h8000149C: output_data <= 32'b10101111111000100000000001111000;
                            32'h800014A0: output_data <= 32'b10101111111111010000000001111100;
                            32'h800014A4: output_data <= 32'b10001111111000010000000000000000;
                            32'h800014A8: output_data <= 32'b10001111111000100000000000000100;
                            32'h800014AC: output_data <= 32'b10001111111000110000000000001000;
                            32'h800014B0: output_data <= 32'b10001111111001000000000000001100;
                            32'h800014B4: output_data <= 32'b10001111111001010000000000010000;
                            32'h800014B8: output_data <= 32'b10001111111001100000000000010100;
                            32'h800014BC: output_data <= 32'b10001111111001110000000000011000;
                            32'h800014C0: output_data <= 32'b10001111111010000000000000011100;
                            32'h800014C4: output_data <= 32'b10001111111010010000000000100000;
                            32'h800014C8: output_data <= 32'b10001111111010100000000000100100;
                            32'h800014CC: output_data <= 32'b10001111111010110000000000101000;
                            32'h800014D0: output_data <= 32'b10001111111011000000000000101100;
                            32'h800014D4: output_data <= 32'b10001111111011010000000000110000;
                            32'h800014D8: output_data <= 32'b10001111111011100000000000110100;
                            32'h800014DC: output_data <= 32'b10001111111011110000000000111000;
                            32'h800014E0: output_data <= 32'b10001111111100000000000000111100;
                            32'h800014E4: output_data <= 32'b10001111111100010000000001000000;
                            32'h800014E8: output_data <= 32'b10001111111100100000000001000100;
                            32'h800014EC: output_data <= 32'b10001111111100110000000001001000;
                            32'h800014F0: output_data <= 32'b10001111111101000000000001001100;
                            32'h800014F4: output_data <= 32'b10001111111101010000000001010000;
                            32'h800014F8: output_data <= 32'b10001111111101100000000001010100;
                            32'h800014FC: output_data <= 32'b10001111111101110000000001011000;
                            32'h80001500: output_data <= 32'b10001111111110000000000001011100;
                            32'h80001504: output_data <= 32'b10001111111110010000000001100000;
                            32'h80001508: output_data <= 32'b10001111111111000000000001101100;
                            32'h8000150C: output_data <= 32'b10001111111111010000000001110000;
                            32'h80001510: output_data <= 32'b10001111111111100000000001110100;
                            32'h80001514: output_data <= 32'b00111100000111111000000000000000;
                            32'h80001518: output_data <= 32'b00100111111111110001010100101000;
                            32'h80001520: output_data <= 32'b00000011010000000000000000001000;
                            32'h8000152C: output_data <= 32'b00111100000111111000000001111111;
                            32'h80001530: output_data <= 32'b00100111111111110000000000000000;
                            32'h80001534: output_data <= 32'b10101111111000010000000000000000;
                            32'h80001538: output_data <= 32'b10101111111000100000000000000100;
                            32'h8000153C: output_data <= 32'b10101111111000110000000000001000;
                            32'h80001540: output_data <= 32'b10101111111001000000000000001100;
                            32'h80001544: output_data <= 32'b10101111111001010000000000010000;
                            32'h80001548: output_data <= 32'b10101111111001100000000000010100;
                            32'h8000154C: output_data <= 32'b10101111111001110000000000011000;
                            32'h80001550: output_data <= 32'b10101111111010000000000000011100;
                            32'h80001554: output_data <= 32'b10101111111010010000000000100000;
                            32'h80001558: output_data <= 32'b10101111111010100000000000100100;
                            32'h8000155C: output_data <= 32'b10101111111010110000000000101000;
                            32'h80001560: output_data <= 32'b10101111111011000000000000101100;
                            32'h80001564: output_data <= 32'b10101111111011010000000000110000;
                            32'h80001568: output_data <= 32'b10101111111011100000000000110100;
                            32'h8000156C: output_data <= 32'b10101111111011110000000000111000;
                            32'h80001570: output_data <= 32'b10101111111100000000000000111100;
                            32'h80001574: output_data <= 32'b10101111111100010000000001000000;
                            32'h80001578: output_data <= 32'b10101111111100100000000001000100;
                            32'h8000157C: output_data <= 32'b10101111111100110000000001001000;
                            32'h80001580: output_data <= 32'b10101111111101000000000001001100;
                            32'h80001584: output_data <= 32'b10101111111101010000000001010000;
                            32'h80001588: output_data <= 32'b10101111111101100000000001010100;
                            32'h8000158C: output_data <= 32'b10101111111101110000000001011000;
                            32'h80001590: output_data <= 32'b10101111111110000000000001011100;
                            32'h80001594: output_data <= 32'b10101111111110010000000001100000;
                            32'h80001598: output_data <= 32'b10101111111111000000000001101100;
                            32'h8000159C: output_data <= 32'b10101111111111010000000001110000;
                            32'h800015A0: output_data <= 32'b10101111111111100000000001110100;
                            32'h800015A4: output_data <= 32'b10001111111111010000000001111100;
                            32'h800015A8: output_data <= 32'b00110100000001000000000000000111;
                            32'h800015AC: output_data <= 32'b00001100000000000000010101110011;
                            32'h800015B4: output_data <= 32'b00001000000000000000010101101111;
                            32'h800015BC: output_data <= 32'b00001000000000000000010010111001;
                            32'h800015C4: output_data <= 32'b00010000000000001111111111111111;
                            32'h800015CC: output_data <= 32'b00111100000010011011111111010000;
                            32'h800015D0: output_data <= 32'b10000001001010000000001111111100;
                            32'h800015D4: output_data <= 32'b00110001000010000000000000000001;
                            32'h800015D8: output_data <= 32'b00010101000000000000000000000011;
                            32'h800015E0: output_data <= 32'b00001000000000000000010101110100;
                            32'h800015E8: output_data <= 32'b00111100000010011011111111010000;
                            32'h800015EC: output_data <= 32'b10100001001001000000001111111000;
                            32'h800015F0: output_data <= 32'b00000011111000000000000000001000;
                            32'h800015F8: output_data <= 32'b00111100000010011011111111010000;
                            32'h800015FC: output_data <= 32'b10000001001010000000001111111100;
                            32'h80001600: output_data <= 32'b00110001000010000000000000000010;
                            32'h80001604: output_data <= 32'b00010101000000000000000000000011;
                            32'h8000160C: output_data <= 32'b00001000000000000000010101111111;
                            32'h80001614: output_data <= 32'b00111100000010011011111111010000;
                            32'h80001618: output_data <= 32'b10000001001000100000001111111000;
                            32'h8000161C: output_data <= 32'b00000011111000000000000000001000;
                            32'h80001624: output_data <= 32'b00100111101111011111111111101100;
                            32'h80001628: output_data <= 32'b10101111101111110000000000000000;
                            32'h8000162C: output_data <= 32'b10101111101100000000000000000100;
                            32'h80001630: output_data <= 32'b10101111101100010000000000001000;
                            32'h80001634: output_data <= 32'b10101111101100100000000000001100;
                            32'h80001638: output_data <= 32'b10101111101100110000000000010000;
                            32'h8000163C: output_data <= 32'b00001100000000000000010101111110;
                            32'h80001644: output_data <= 32'b00000000000000101000000000100101;
                            32'h80001648: output_data <= 32'b00001100000000000000010101111110;
                            32'h80001650: output_data <= 32'b00000000000000101000100000100101;
                            32'h80001654: output_data <= 32'b00001100000000000000010101111110;
                            32'h8000165C: output_data <= 32'b00000000000000101001000000100101;
                            32'h80001660: output_data <= 32'b00001100000000000000010101111110;
                            32'h80001668: output_data <= 32'b00000000000000101001100000100101;
                            32'h8000166C: output_data <= 32'b00110010000100000000000011111111;
                            32'h80001670: output_data <= 32'b00110010011100110000000011111111;
                            32'h80001674: output_data <= 32'b00110010010100100000000011111111;
                            32'h80001678: output_data <= 32'b00110010001100010000000011111111;
                            32'h8000167C: output_data <= 32'b00000000000100110001000000100101;
                            32'h80001680: output_data <= 32'b00000000000000100001001000000000;
                            32'h80001684: output_data <= 32'b00000000010100100001000000100101;
                            32'h80001688: output_data <= 32'b00000000000000100001001000000000;
                            32'h8000168C: output_data <= 32'b00000000010100010001000000100101;
                            32'h80001690: output_data <= 32'b00000000000000100001001000000000;
                            32'h80001694: output_data <= 32'b00000000010100000001000000100101;
                            32'h80001698: output_data <= 32'b10001111101111110000000000000000;
                            32'h8000169C: output_data <= 32'b10001111101100000000000000000100;
                            32'h800016A0: output_data <= 32'b10001111101100010000000000001000;
                            32'h800016A4: output_data <= 32'b10001111101100100000000000001100;
                            32'h800016A8: output_data <= 32'b10001111101100110000000000010000;
                            32'h800016AC: output_data <= 32'b00100111101111010000000000010100;
                            32'h800016B0: output_data <= 32'b00000011111000000000000000001000;
                            default: begin
                                if (addr[31:20]==12'h800)
                                    output_data <= 32'b0;
                                else
                                    output_data <= ram_read_data;
                            end
                        endcase
*/
                        output_data <= ram_read_data;

                        be <= 4'b0000; 
                    end
                end
                else if (if_write) begin
                    if (bytemode) begin
                        case (addr[1:0])
                            2'b00: begin
                                ram_write_data <= {input_data[7:0], 24'b0};
                                be <= 4'b0111;
                            end
                            2'b01: begin
                                ram_write_data <= {8'b0, input_data[7:0], 16'b0};
                                be <= 4'b1011;
                            end
                            2'b10: begin
                                ram_write_data <= {16'b0, input_data[7:0], 8'b0};
                                be <= 4'b1101;
                            end
                            2'b11: begin
                                ram_write_data <= {24'b0, input_data[7:0]};
                                be <= 4'b1110;
                            end
                            default: begin
                                ram_write_data <= input_data;
                                be <= 4'b0000;
                            end
                        endcase
                    end
                    else begin
                        ram_write_data <= input_data;
                        be <= 4'b0000; 
                    end
                end
            end
        endcase
    end
    else begin
        // ram
        ce1 <= 1'b1;
        ce2 <= 1'b1;
        oe1 <= 1'b1;
        oe2 <= 1'b1;
        we1 <= 1'b1;
        we2 <= 1'b1;
        rdn <= 1'b1;
        wrn <= 1'b1;
    end
end

endmodule
